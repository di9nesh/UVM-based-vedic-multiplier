import uvm_pkg::*;
`include "uvm_macros.svh"
import ved_pkg::*;

class ved_test_corner extends ved_base_test;
  `uvm_component_utils(ved_test_corner)

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  task run_phase(uvm_phase phase);
    ved_corner_seq seq;

    phase.raise_objection(this);

    seq = ved_corner_seq::type_id::create("seq");
    seq.start(env.agt.sqr);

    repeat (10) @(posedge env.agt.vif.clk);

    phase.drop_objection(this);
  endtask
endclass

